module org(
  input x, y,
  output z);
  or(z,x,y);
endmodule
