
module xor_gate (A,B,Y);
  input A,B;
  output Y;
  xor(Y,A,B);
endmodule
