module andg(
  input x, y,
  output z);
  and(z,x,y);
endmodule
